module testbench();
reg [31:0] a,b;
reg clk;
wire [31:0] out;

FPU32bitAdderTop test(a,b,clk,out);
initial 
begin 
clk=1'b0;
a=32'b01000000011010011110001101010100; //3.6545
b=32'b01000000101110000111111111001100; //5.7656
#50;
a=32'b01000010110010001110100111011011; //100.45675
b=32'b01000001000111100000011000100101; //9.8765
#50;
a=32'b01000001001100011100011100010001; //11.1111
b=32'b00000000000000000000000000000000; //0
#50;
$stop;
end
always #10 clk=!clk;
endmodule