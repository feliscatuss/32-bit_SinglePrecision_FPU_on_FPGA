`timescale 1ps / 1ps

module FPU32bitAdderTB;

	reg clk;
	reg [31:0] a, b;

	wire [31:0] out;

	FPU32bitAdderTop uut (a, b, clk, out); 

	initial 
	begin
		clk = 0;
		a = 0;
		b = 0;
#10;
      clk = 0;
		a = 32'b11000000100100110011001100110011;//-4.6
		b = 32'b11000000100100110011001100110011;//-4.6
		//out = 11000001000100110011001100110011;//-9.2
#20;
		clk = 0;
		a = 32'b11000000100100110011001100110011;//-4.6;
		b = 32'b00111111000110011001100110011001;//0.6
		//out = 11000000100000000000000000000000 //-4
#30;
    	clk = 0;
		a = 32'b01000000010011001100110011001100;//3.2;
		b = 32'b10111111000110011001100110011001;//-0.6
		//out = 01000000001001100110011001100110 //2.6

#40;
 	   clk = 0;
		a = 32'b01000101000010100111000011001100;//2215.05;
		b = 32'b01000101000010011101000110011001;//2205.10
		//out = 01000101100010100010000100110011 //4420.15

#50;
   end	
   always #5 clk=(~clk);  
endmodule